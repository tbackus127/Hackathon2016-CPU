module jump (offset);

input [15:0]offset;


end module


module jump_less_than(ComparatorA, ComapatorB, offset);

input [15:0]ComparatorA;
input [15:0]ComparatorB;
input [4:0]offset;

if (ComparatorA[15] < ComparatorB[15])
    
if (ComparatorA[14] < ComparatorB[14])

if (ComparatorA[13] < ComparatorB[13])

if (ComparatorA[12] < ComparatorB[12])

if (ComparatorA[11] < ComparatorB[11])

if (ComparatorA[10] < ComparatorB[10])

if (ComparatorA[9] < ComparatorB[9])

if (ComparatorA[8] < ComparatorB[8])

if (ComparatorA[7] < ComparatorB[7])

if (ComparatorA[6] < ComparatorB[6])

if (ComparatorA[5] < ComparatorB[5])

if (ComparatorA[4] < ComparatorB[4])

if (ComparatorA[3] < ComparatorB[3])

if (ComparatorA[2] < ComparatorB[2])

if (ComparatorA[1] < ComparatorB[1])

if (ComparatorA[0] < ComparatorB[0]);

end module
