module program_counter (regOP, newReg, offset);

input [15:0]regOP;
output [15:0]newReg;

assign newReg[0] = ;
assign newReg[1] = ;
assign newReg[2] = ;
assign newReg[3] = ;
assign newReg[4] = ;
assign newReg[5] = ;
assign newReg[6] = ;
assign newReg[7] = ;
assign newReg[8] = ;
assign newReg[9] = ;
assign newReg[10] = ;
assign newReg[11] = ;
assign newReg[12] = ;
assign newReg[13] = ;
assign newReg[14] = ;
assign newReg[15] = ;

end module
